// Diseño:      rom_mul
// Archivo:     rom_mul_tb.v
// Descripción: Multiplicador basado en ROM
// Autor:       Jorge Juan <jjchico@gmail.com>
// Fecha:       11/06/2010

/*
   Lección 8-1. Multiplicador basado en ROM.

   Este archivo contiene un banco de pruebas para verificar las diferentes
   operaciones del multiplicador basado en ROM en rom_mul.v.
*/

`timescale 1ns / 1ps

// Banco de pruebas

module test();

endmodule // test


/*
   EJERCICIOS

*/
